class Agent

endclass
