class Agent extends  /* base class*/;
	
endclass : Agent